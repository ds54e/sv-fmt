module comment_demo;
  initial begin

    /*block*/

    assign a = 1; //inline
  end
endmodule
