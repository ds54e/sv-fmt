module randseq_demo;
initial begin
randsequence(req)
req : { foo = 1; };
endsequence
end
endmodule
