module randcase_demo;
initial begin
randcase
  10: data <= 1;
  1: data <= 0;
endcase
end
endmodule
